module ALU{
	.data1_i,
	.data2_i,
	.ALUControl_i,
	.data_o
};

//Ports
