module ID_EX(
	clk_i,
	WB_i,
	WB_o,
	M_i,
	M_o,
	EX_i,
	EX_o_1,
	EX_o_2,
	EX_o_3,
	PC_i,
	ReadData1_i,	//RS
	ReadData2_i,	//RT
	inst1_i,
	inst2_i,
	inst3_i,
	inst4_i,
	inst5_i,
	MUX6_o,
	MUX7_o,
	inst1_o,	//MUX4_o
	inst2_o,
	inst3_o,
	inst4_o,
	inst5_o,
	stall
);

input clk_i, stall;
input   [3:0]   EX_i;
input   [1:0]WB_i;
input	[2:0]M_i;
input 	[31:0]	PC_i;
input   [31:0]ReadData1_i, ReadData2_i;
output  reg [1:0]WB_o;
output  reg [2:0]M_o;
output  reg EX_o_1, EX_o_3;
output  reg [1:0]EX_o_2;
input	[31:0]	inst1_i;
input   [4:0]	inst2_i, inst3_i, inst4_i, inst5_i;
output	reg [31:0]inst1_o;
output  reg [4:0]inst2_o, inst3_o, inst4_o, inst5_o;
output  reg [31:0]MUX6_o, MUX7_o;


always @(posedge clk_i) begin
	if(stall == 1'b1) begin
		
	end
	else begin
    WB_o = WB_i;
    M_o = M_i;
    //TODO EX!!
    EX_o_1 = EX_i[3];
    EX_o_2 = EX_i[2:1];
    EX_o_3 = EX_i[0];
    inst1_o = inst1_i;
    inst2_o = inst2_i;
    inst3_o = inst3_i;
    inst4_o = inst4_i;
    inst5_o = inst5_i;
    MUX6_o  = ReadData1_i;
    MUX7_o  = ReadData2_i;
	end
end

endmodule


